pll_inst : pll PORT MAP (
		inclk0	 => inclk0_sig,	-- in
		c0	 => c0_sig					-- out
	);

